library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity name is
    generic 
    (

    );
    port 
    (

    );
end entity;

architecture behavorial of name is
    signal
begin

end architecture;
